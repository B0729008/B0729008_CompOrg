// Copyright (C) 1991-2010 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II"
// VERSION		"Version 10.0 Build 218 06/27/2010 SJ Web Edition"
// CREATED		"Fri Oct 25 16:24:24 2019"

module Block2(
	S1,
	A,
	B,
	C,
	D,
	S0,
	Q
);


input wire	S1;
input wire	A;
input wire	B;
input wire	C;
input wire	D;
input wire	S0;
output wire	Q;

wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;




assign	SYNTHESIZED_WIRE_4 = S1 & S0 & A;

assign	SYNTHESIZED_WIRE_7 = S1 & SYNTHESIZED_WIRE_8 & B;

assign	SYNTHESIZED_WIRE_5 = SYNTHESIZED_WIRE_9 & S0 & C;

assign	SYNTHESIZED_WIRE_6 = SYNTHESIZED_WIRE_9 & SYNTHESIZED_WIRE_8 & D;

assign	Q = SYNTHESIZED_WIRE_4 | SYNTHESIZED_WIRE_5 | SYNTHESIZED_WIRE_6 | SYNTHESIZED_WIRE_7;

assign	SYNTHESIZED_WIRE_9 =  ~S1;

assign	SYNTHESIZED_WIRE_8 =  ~S0;


endmodule
