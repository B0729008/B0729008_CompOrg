library verilog;
use verilog.vl_types.all;
entity lab05 is
    port(
        clk             : in     vl_logic;
        clean           : in     vl_logic;
        lout0a          : out    vl_logic;
        lout0b          : out    vl_logic;
        lout0c          : out    vl_logic;
        lout0d          : out    vl_logic;
        lout0e          : out    vl_logic;
        lout0f          : out    vl_logic;
        lout0g          : out    vl_logic;
        lout1a          : out    vl_logic;
        lout1b          : out    vl_logic;
        lout1c          : out    vl_logic;
        lout1d          : out    vl_logic;
        lout1e          : out    vl_logic;
        lout1f          : out    vl_logic;
        lout1g          : out    vl_logic;
        lout2a          : out    vl_logic;
        lout2b          : out    vl_logic;
        lout2c          : out    vl_logic;
        lout2d          : out    vl_logic;
        lout2e          : out    vl_logic;
        lout2f          : out    vl_logic;
        lout2g          : out    vl_logic;
        lout3a          : out    vl_logic;
        lout3b          : out    vl_logic;
        lout3c          : out    vl_logic;
        lout3d          : out    vl_logic;
        lout3e          : out    vl_logic;
        lout3f          : out    vl_logic;
        lout3g          : out    vl_logic
    );
end lab05;
